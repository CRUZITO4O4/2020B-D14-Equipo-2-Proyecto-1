module sumador2(
	input[31:0]inputsumador1,inputsumador2,
	output[31:0]outputsumador
);

assign outputsumador = inputsumador1 + inputsumador2;

endmodule
