module Comp_AND(
	input inputand1,
	input inputand2,
	output outputand
);

assign outputand = inputand1 & inputand2;

endmodule
